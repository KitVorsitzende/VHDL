library verilog;
use verilog.vl_types.all;
entity Faltungscodierer_vlg_vec_tst is
end Faltungscodierer_vlg_vec_tst;
